//Subject:     CO project 2 - Decoder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      Luke,0816192
//----------------------------------------------
//Date:        2010/8/16
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Decoder(
    instr_op_i,
	RegWrite_o,
	ALU_op_o,
	ALUSrc_o,
	RegDst_o,
	Branch_o,
	Jump_o,
	MemRead_o,
	MemWrite_o,
	MemtoReg_o
	);
     
//I/O ports
input  [6-1:0] instr_op_i;

output         RegWrite_o;
output [3-1:0] ALU_op_o;
output         ALUSrc_o;
output [2-1:0] RegDst_o;
output         Branch_o;
output 		   Jump_o;
output		   MemRead_o;
output		   MemWrite_o;
output [2-1:0] MemtoReg_o;
 
//Internal Signals
reg    [3-1:0] ALU_op_o;
reg            ALUSrc_o;
reg            RegWrite_o;
reg	   [2-1:0] RegDst_o;
reg            Branch_o;
reg 		      Jump_o;
reg			   MemRead_o;
reg			   MemWrite_o;
reg	   [2-1:0] MemtoReg_o;

wire		   R_ctrl;
wire		   lw_ctrl;
wire		   sw_ctrl;
wire		   beq_ctrl;
wire		   addi_ctrl;
wire		   slti_ctrl;
wire		   j_ctrl;
wire		   jal_ctrl;


assign R_ctrl = &(~instr_op_i);

assign lw_ctrl	= (instr_op_i== 6'b100011);
assign sw_ctrl	= (instr_op_i== 6'b101011);
assign beq_ctrl	= (instr_op_i== 6'd4);
assign addi_ctrl	= (instr_op_i== 6'd8);
assign slti_ctrl	= (instr_op_i== 6'd10);

assign j_ctrl	= (instr_op_i== 6'b000010);
assign jal_ctrl	= (instr_op_i== 6'b000011);

always @(instr_op_i)begin
    Branch_o <= beq_ctrl;
    
    if(lw_ctrl)
		MemtoReg_o <= 1;
	else if(jal_ctrl)
		MemtoReg_o <= 2;
	else
		MemtoReg_o <= 0;
	
	Jump_o <= j_ctrl | jal_ctrl;
	MemRead_o <= lw_ctrl;
	MemWrite_o <= sw_ctrl;	
	ALUSrc_o <= addi_ctrl | slti_ctrl | lw_ctrl | sw_ctrl;
	RegWrite_o <= R_ctrl | addi_ctrl | slti_ctrl | lw_ctrl | jal_ctrl;
	RegDst_o <= R_ctrl ? 1:(jal_ctrl ? 2 : 0);
end

always @(instr_op_i)begin
	if(lw_ctrl | sw_ctrl)
		ALU_op_o <= 3'd0; // lw or sw
	else if(beq_ctrl)
		ALU_op_o <= 3'd1; // beq
	else if(R_ctrl)
		ALU_op_o <= 3'd2; // R
	else if(addi_ctrl)
		ALU_op_o <= 3'd3; // 3 addi
	else if(slti_ctrl)
		ALU_op_o <= 3'd4; // 4 slti
	else
		ALU_op_o <= 3'b111;
end

endmodule





                    
                    